// ECE 5440: Advanced Digital Design
// Author: Matthew Andersen 2071
// RNG_LFSR_3b
// This takes an enable signal and outputs
// a random 3-bit number. The number is pseudo random b/c
// 50 MHz clock means any random time interval between getting the numbers
// results in a random 3 bit output.

module RNG_LFSR_3b(RNG_Gen, Random_Num, clk, rst);
   input RNG_Gen, clk, rst;
   output [2:0] Random_Num;
   reg [15:0] LFSR;
   wire feedback = LFSR[15];
   
   assign Random_Num = {LFSR[1], LFSR[5], LFSR[10]};

   always @(posedge clk)
   begin
      if (rst == 1'b0) begin
        LFSR <= 16'b0000000000000000;
      end
      else begin
         if (RNG_Gen == 1'b1) begin
            LFSR[0] <= feedback;
            LFSR[1] <= LFSR[0];
            LFSR[2] <= LFSR[1] ~^ feedback;
            LFSR[3] <= LFSR[2] ~^ feedback;
            LFSR[4] <= LFSR[3];
            LFSR[5] <= LFSR[4] ~^ feedback;
            LFSR[6] <= LFSR[5];
            LFSR[7] <= LFSR[6];
            LFSR[8] <= LFSR[7];
            LFSR[9] <= LFSR[8];
            LFSR[10] <= LFSR[9];
            LFSR[11] <= LFSR[10];
            LFSR[12] <= LFSR[11];
            LFSR[13] <= LFSR[12];
            LFSR[14] <= LFSR[13];
            LFSR[15] <= LFSR[14];
         end
      end
   end
endmodule